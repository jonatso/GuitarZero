`ifndef __TINY_SYNTH_TONE_TRIANGLE__
`define __TINY_SYNTH_TONE_TRIANGLE__
/* =============================
 * Triangle tone generator
 * =============================
 *
 * Generates a triangle-wave; optionally ring-modulated with the MSB of
 * another oscillator.
 *
 * Principle of operation:
 *
 * Since we want the triangle wave to count up, and back down while the
 * accumulator transitions from 0 to full-scale, we need a way of inverting
 * the wave at half-scale.
 *
 * It turns out that binary inverting a counter makes it count in the
 * reverse direction, so we use the accumulator MSB to optionally invert
 * the bottom bits of the accumulator, which are then shifted into the
 * output.
 *
 * The "inversion" of the counter can also be driven by the MSB
 * from another oscillator, and in SID terms this is known as "ring modulation".
 * This allows for some quite complex waveforms to be generated by connecting
 * multiple voices together.
 */
module tone_generator_triangle #(
  parameter ACCUMULATOR_BITS = 24,
  parameter OUTPUT_BITS = 12)
(
  input [ACCUMULATOR_BITS-1:0] accumulator,
  output wire [OUTPUT_BITS-1:0] dout);

  wire invert_wave;

  // invert the waveform (ie. start counting down instead of up)
  // if either ringmod is enabled and high,
  // or MSB of accumulator is set.
  assign invert_wave = accumulator[ACCUMULATOR_BITS-1];

  assign dout = invert_wave ? ~accumulator[ACCUMULATOR_BITS-2 -: OUTPUT_BITS]
                            : accumulator[ACCUMULATOR_BITS-2 -: OUTPUT_BITS];

endmodule

`endif
